library IEEE;
use IEEE.std_logic_1164.ALL;
use IEEE.numeric_std.ALL;


entity rom256x16 is
  port (
    clk: in std_logic;
    A: in std_logic_vector(8-1 downto 0);
    D: out std_logic_vector(16-1 downto 0)
  );
end entity rom256x16;


architecture behav of rom256x16 is
begin
  process (clk)
  begin
    if rising_edge(clk) then
       case A is

---   when x"00" => D <= "0111000001101110";
---   when x"01" => D <= "1001000000000000";
---   when x"02" => D <= "1000000000000000";
---   when x"03" => D <= "0111001000010100";
---   when x"04" => D <= "0111010001100100";
---   when x"05" => D <= "0111110000000010";
---   when x"06" => D <= "0001010010011010";
---   when x"07" => D <= "0001011000011001";
---   when x"08" => D <= "0001011110011011";
---   when x"09" => D <= "0001011010011011";
---   when x"0a" => D <= "0001010011010001";
---   when x"0b" => D <= "1001010000000001";
---   when x"0c" => D <= "0011001001000001";
---   when x"0d" => D <= "1110000000001111";
---   when x"0e" => D <= "1111000000000110";
---   when others => D <= x"0000";

---when x"00" => D <= "0111000000100000";
---when x"01" => D <= "1001000000000001";
---when x"02" => D <= "1000001000000001";
---when x"03" => D <= "0111010001100100";
---when x"04" => D <= "0111101000000010";
---when x"05" => D <= "0111110000001010";
---when x"06" => D <= "0001010010011010";
---when x"07" => D <= "0001011001011000";
---when x"08" => D <= "0001011101011011";
---when x"09" => D <= "0001011010010011";
---when x"0a" => D <= "0011110110000001";
---when x"0b" => D <= "1110000000001101";
---when x"0c" => D <= "1111000000000110";
---when x"0d" => D <= "1001010000000001";
---when others => D <= x"0000";
---
when x"00" => D <= "0111000000001010";
when x"01" => D <= "1001000000000000";
when x"02" => D <= "1000000000000000";
when x"03" => D <= "0111001000010110";
when x"04" => D <= "0111010000000111";
when x"05" => D <= "0001000000000010";
when x"06" => D <= "0001000001000010";
when x"07" => D <= "0001000010000011";
when x"08" => D <= "1001000000000001";
when others => D <= x"0000";



       end case; 
    end if;
  end process;
end behav;
